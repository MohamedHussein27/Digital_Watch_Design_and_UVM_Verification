package dw_agent_pkg;
    import dw_config_obj_pkg::*;
    import dw_driver_pkg::*;
    import dw_monitor_pkg::*;
    import dw_seq_item_pkg::*;
    import dw_sequencer_pkg::*;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    class dw_agent extends uvm_agent;
        `uvm_component_utils(dw_agent)

        dw_config_obj dw_cfg; // configuration object
        dw_driver drv; // driver
        dw_monitor mon; // monitor
        dw_sequencer sqr; // sequencer
        
        uvm_analysis_port #(dw_seq_item) agt_ap; // will be used to connect scoreboard and coverage collector

        function new (string name = "dw_agent", uvm_component parent = null);
            super.new(name, parent);
        endfunction

        function void build_phase(uvm_phase phase);
            super.build_phase(phase);
            if(!uvm_config_db #(dw_config_obj)::get(this,"","CFG", dw_cfg)) begin
                    `uvm_fatal("build_phase","agent error");
            end
            // creation
            drv = dw_driver::type_id::create("driver", this);
            mon = dw_monitor::type_id::create("mon", this);
            sqr = dw_sequencer::type_id::create("sqr", this);
            agt_ap = new("agt_ap", this); // connection point
        endfunction

        function void connect_phase(uvm_phase phase);
            super.connect_phase(phase);
            drv.dw_vif = dw_cfg.dw_vif;
            mon.dw_vif = dw_cfg.dw_vif;
            drv.seq_item_port.connect(sqr.seq_item_export);
            mon.mon_ap.connect(agt_ap); // connect monitor share point with agent share point so the monitor will be able to get data from the scoreboard and the cov collector
        endfunction
    endclass
endpackage